module bpl2a(chaves,t1,t2);
	input [7:0] chaves;
	output [6:0] t1,t2;
	
endmodule 