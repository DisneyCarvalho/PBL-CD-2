module ejdjds(A,S);
	input [5:0] A;
	output [5:0] S;
	
	not(S,A);
	
	
endmodule 