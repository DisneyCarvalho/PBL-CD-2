module fafafgga(a,b,s);
	input a,b;
	output [3:0] s;
	
	wire fio1;
	
	somadorcompleto(a,b,0,s,fio1);
	
endmodule 

