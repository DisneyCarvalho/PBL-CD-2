module bpl2 (clock,l1,c1);
	input [18:0] clock;
	output l1,c1;
	
	
	
	always @(posedge clock) begin 
	
	end
	
	
endmodule 